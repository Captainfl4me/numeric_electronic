-------------------------------------------------------
-- Ce programme a été développé à CENTRALE-SUPELEC
-- Merci de conserver ce cartouche
-- Copyright  (c) 2022  CENTRALE-SUPELEC   
-- Département Systèmes électroniques
-- ---------------------------------------------------
--
-- fichier : testbench_e.vhd
-- auteur  : P.BENABES   
-- Copyright (c) 2022 CENTRALE-SUPELEC
-- Revision: 4.1  Date: 22/02/2022
--
-- ---------------------------------------------------
-- ---------------------------------------------------
--
-- DESCRIPTION DU SCRIPT :
-- entité du testbench
--
--------------------------------------------------------

library IEEE;
use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.fixed_float_types.all;	-- package virgule fixe
use ieee.fixed_pkg.all;
use ieee.math_real.all;			-- bibliotheque mathématique pour la trigonométrie
use work.types.all ;			-- les types predefinis

entity testbench  is
end testbench;


